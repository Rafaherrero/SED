--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   17:00:06 02/23/2014
-- Design Name:   
-- Module Name:   C:/Users/Rafa/practica/funciones_tb.vhd
-- Project Name:  practica
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: funciones
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY funciones_tb IS
END funciones_tb;
 
ARCHITECTURE behavior OF funciones_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT funciones
    PORT(
         a : IN  std_logic;
         b : IN  std_logic;
         fnot : OUT  std_logic;
         fand : OUT  std_logic;
         ffor : OUT  std_logic;
         fnand : OUT  std_logic;
         fnor : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal a : std_logic := '0';
   signal b : std_logic := '0';

 	--Outputs
   signal fnot : std_logic;
   signal fand : std_logic;
   signal ffor : std_logic;
   signal fnand : std_logic;
   signal fnor : std_logic;
  
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: funciones PORT MAP (
          a => a,
          b => b,
          fnot => fnot,
          fand => fand,
          ffor => ffor,
          fnand => fnand,
          fnor => fnor
        );
		  
		  a <= not a after 10 ns;
		  b <= not b after 20 ns;
END;
