--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   23:33:36 05/11/2014
-- Design Name:   
-- Module Name:   C:/Users/Rafa/Desktop/probando/pfinal/pfinal/cronometro_tb.vhd
-- Project Name:  pfinal
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: cronometro
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY cronometro_tb IS
END cronometro_tb;
 
ARCHITECTURE behavior OF cronometro_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT cronometro
    PORT(
         clk : IN  std_logic;
         reset : IN  std_logic;
         ce : IN  std_logic;
         botons : IN  std_logic;
         botonm : IN  std_logic;
         ledce : IN  std_logic;
         sd : OUT  std_logic_vector(6 downto 0);
         an0 : OUT  std_logic;
         an1 : OUT  std_logic;
         an2 : OUT  std_logic;
         an3 : OUT  std_logic;
         ledsalida : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal reset : std_logic := '0';
   signal ce : std_logic := '0';
   signal botons : std_logic := '0';
   signal botonm : std_logic := '0';
   signal ledce : std_logic := '0';

 	--Outputs
   signal sd : std_logic_vector(6 downto 0);
   signal an0 : std_logic;
   signal an1 : std_logic;
   signal an2 : std_logic;
   signal an3 : std_logic;
   signal ledsalida : std_logic;

   -- Clock period definitions
   constant clk_period : time := 20 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: cronometro PORT MAP (
          clk => clk,
          reset => reset,
          ce => ce,
          botons => botons,
          botonm => botonm,
          ledce => ledce,
          sd => sd,
          an0 => an0,
          an1 => an1,
          an2 => an2,
          an3 => an3,
          ledsalida => ledsalida
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      wait for clk_period*10;

      -- insert stimulus here 

      wait;
   end process;

END;
